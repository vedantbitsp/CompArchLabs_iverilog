module 4bit_comparator (a , b, , x , y, z);
input [3:0]a, [3:0]b;
output x, y, z;

